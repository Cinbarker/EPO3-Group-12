library IEEE;
use IEEE.std_logic_1164.ALL;

entity clearing3_tb is
end clearing3_tb;

