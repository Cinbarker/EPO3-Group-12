configuration controller_fsm_tb_behaviour_tb_cfg of controller_fsm_tb is
   for behaviour_tb
      for all: controller_fsm use configuration work.controller_fsm_behaviour_cfg;
      end for;
   end for;
end controller_fsm_tb_behaviour_tb_cfg;
