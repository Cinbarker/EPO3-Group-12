library IEEE;
use IEEE.std_logic_1164.ALL;

entity pulse_gen_tb is
end pulse_gen_tb;

