configuration clearing3_behaviour_cfg of clearing3 is
   for behaviour
   end for;
end clearing3_behaviour_cfg;
