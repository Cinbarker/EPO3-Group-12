library IEEE;
use IEEE.std_logic_1164.ALL;

entity minecounter_tb is
end minecounter_tb;

