configuration controller_fsm_behaviour_cfg of controller_fsm is
   for behaviour
   end for;
end controller_fsm_behaviour_cfg;
