library IEEE;
use IEEE.std_logic_1164.ALL;

entity seedgen_tb is
end seedgen_tb;

