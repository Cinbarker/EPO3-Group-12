library IEEE;
use IEEE.std_logic_1164.ALL;

entity controller_fsm_tb is
end controller_fsm_tb;

