library IEEE;
use IEEE.std_logic_1164.ALL;  
use IEEE.numeric_std.ALL;
entity maps is

   port(x_address : in  std_logic_vector(3 downto 0);
	y_address : in  std_logic_vector(3 downto 0);

        data    : out std_logic_vector(5 downto 0));	--red(1)red(0)green(1)green(0)blue(1)b1ue(0) (rrggbb)

end maps;  

library IEEE;

use IEEE.std_logic_1164.ALL;  

architecture behaviour of rom is

type bitmap is array (0 to 10, 0 to 10) of std_logic_vector (5 downto 0);			-- this creates an 11 by 11 matrix see below
signal mine_map : bitmap := (	("111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111"),
				("111111", "111111", "111111", "111111", "111111", "000000", "111111", "111111", "111111", "111111", "111111"),
				("111111", "111111", "000000", "111111", "111111", "000000", "111111", "111111", "000000", "111111", "111111"),
				("111111", "111111", "111111", "000000", "000000", "000000", "000000", "000000", "111111", "111111", "111111"),
				("111111", "111111", "111111", "000000", "111111", "000000", "000000", "000000", "111111", "111111", "111111"),
				("111111", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "111111"),
				("111111", "111111", "111111", "000000", "000000", "000000", "000000", "000000", "111111", "111111", "111111"),
				("111111", "111111", "111111", "000000", "000000", "000000", "000000", "000000", "111111", "111111", "111111"),
				("111111", "111111", "000000", "111111", "111111", "000000", "111111", "111111", "000000", "111111", "111111"),
				("111111", "111111", "111111", "111111", "111111", "000000", "111111", "111111", "111111", "111111", "111111"),
				("111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111"));
begin


	data <= mine_map(to_integer(unsigned(y_address)), to_integer(unsigned(x_address)));		-- y is for columns, x is for rows

end behaviour;
