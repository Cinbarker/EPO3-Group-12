library IEEE;
use IEEE.std_logic_1164.ALL;

entity buildingmodule_tb is
end buildingmodule_tb;

