library IEEE;
use IEEE.std_logic_1164.ALL;

entity mineplacerv2_tb is
end mineplacerv2_tb;

